
 `timescale     10 ps/ 10 ps  
 `define          DELAY 10  

 module     tb_fifo_mem;  

 parameter     ENDTIME      = 40000;  
 
 // DUT Input regs  
 reg     clk;  
 reg     rst_n;  
 reg     write;  
 reg     read;  
 reg     [7:0] data_in;  
 
 // DUT Output wires  
 wire     [7:0] data_out;  
 wire     is_empty;  
 wire     is_full;  
 wire     threshold;  
 wire     overflow;  
 wire     underflow;  
 integer i;  
 
 // DUT Instantiation
 
 fifo_mem tb1 (
   // Outputs  
   data_out, is_full, is_empty, threshold, overflow,   
   underflow,   
   // Inputs  
   clk, rst_n, write, read, data_in  
   );  
   
 // Initial Conditions 

 initial  
      begin  
           clk     = 1'b0;  
           rst_n     = 1'b0;  
           write     = 1'b0;  
           read     = 1'b0;  
           data_in     = 8'd0;  
      end  
      
 // Generating Test Vectors  
 
 initial  
      begin  
           main;  
      end 
      
 task main;  
      fork  
           clock_generator;  
           reset_generator;  
           operation_process;  
           debug_fifo;  
           endsimulation;  
      join  
 endtask  
 
 // clock_generator Task
 task clock_generator;  
      begin  
           forever #`DELAY clk = !clk;  
      end  
 endtask  
 
 // reset_generator Task
 task reset_generator;  
      begin  
           #(`DELAY*2)  
           rst_n = 1'b1;  
           # 7.9  
           rst_n = 1'b0;  
           # 7.09  
           rst_n = 1'b1;  
      end  
 endtask  
 
 //  operation_process task
 task operation_process;  
      begin  
           for (i = 0; i < 17; i = i + 1) begin: WRE  
                #(`DELAY*5)  
                write = 1'b1;  
                data_in = data_in + 8'd1;  
                #(`DELAY*2)  
                write = 1'b0;  
           end  
           #(`DELAY)  
           for (i = 0; i < 17; i = i + 1) begin: RDE  
                #(`DELAY*2)  
                read = 1'b1;  
                #(`DELAY*2)  
                read = 1'b0;  
           end  
      end  
 endtask  
 
 // Debug prints fifo
 task debug_fifo;  
      begin  
           $display("----------------------------------------------");  
           $display("------------------   -----------------------");  
           $display("----------- SIMULATION RESULT ----------------");  
           $display("--------------       -------------------");  
           $display("----------------     ---------------------");  
           $display("----------------------------------------------");  
           $monitor("TIME = %d, write = %b, read = %b, data_in = %h",$time, write, read, data_in);  
      end  
 endtask  
 
 // Self-Checking  
 reg [5:0] waddr, raddr;  
 reg [7:0] mem[64:0];  
 always @ (posedge clk) begin  
      if (~rst_n) begin  
           waddr     <= 6'd0;  
      end  
      else if (write) begin  
           mem[waddr] <= data_in;  
           waddr <= waddr + 1;  
      end  
      $display("TIME = %d, data_out = %d, mem = %d",$time, data_out,mem[raddr]);  
      if (~rst_n) raddr     <= 6'd0;  
      else if (read & (~is_empty)) raddr <= raddr + 1;  
      if (read & (~is_empty)) begin  
           if (mem[raddr]  
            == data_out) begin  
                $display("=== PASS ===== PASS ==== PASS ==== PASS ===");  
                if (raddr == 16) $finish;  
           end  
           else begin  
                $display ("=== FAIL ==== FAIL ==== FAIL ==== FAIL ===");  
                $display("-------------- THE SIMUALTION FINISHED ------------");  
                $finish;  
           end  
      end  
 end  
 
 // endsimulation task
 task endsimulation;  
      begin  
           #ENDTIME  
           $display("-------------- THE SIMULATION FINISHED ------------");  
           $finish;  
      end  
 endtask  
 
 endmodule